000007970C8000EF
0E8000EF12878793
00A3031380001337
FE038EE300034383
11C7879300000797
2BC003130CC000EF
00138393000073B3
800011B7FE731EE3
0120059308018193
0FF0000F02018023
0061802304100313
001003130FF0000F
0FF0000F00618C23
0261802300100313
00B005130FF0000F
00000513030000EF
024000EF028000EF
00F2F2930045D293
084000EF03028293
0302829300F5F293
0000006F078000EF
0FF0000F00A18823
0FF0000F0081C303
FE031AE300137313
000080670101C583
08000E1380002737
01B00E9301C70623
00300E1301D70023
08700E1301C70623
0007022301C70423
0007828300008067
020FFF9301470F83
00570023FE0F8CE3
0007828300178793
00008067FE0294E3
020FFF9301470F83
00570023FE0F8CE3
6563634100008067
2E2E74736554206C
204D4152000A0D2E
000000000A0D4B4F
0000000000000000
